
module progmem (
    // Closk & reset
    input wire clk,
    input wire rstn,

    // PicoRV32 bus interface
    input  wire        valid,
    output wire        ready,
    input  wire [31:0] addr,
    output wire [31:0] rdata
);

  // ============================================================================

  localparam MEM_SIZE_BITS = 10;  // In 32-bit words
  localparam MEM_SIZE = 1 << MEM_SIZE_BITS;
  localparam MEM_ADDR_MASK = 32'h0010_0000;

  // ============================================================================

  wire [MEM_SIZE_BITS-1:0] mem_addr;
  reg  [             31:0] mem_data;
  reg  [             31:0] mem      [0:MEM_SIZE];

  initial begin
    mem['h0000] <= 32'h00000093;
    mem['h0001] <= 32'h00000193;
    mem['h0002] <= 32'h00000213;
    mem['h0003] <= 32'h00000293;
    mem['h0004] <= 32'h00000313;
    mem['h0005] <= 32'h00000393;
    mem['h0006] <= 32'h00000413;
    mem['h0007] <= 32'h00000493;
    mem['h0008] <= 32'h00000513;
    mem['h0009] <= 32'h00000593;
    mem['h000A] <= 32'h00000613;
    mem['h000B] <= 32'h00000693;
    mem['h000C] <= 32'h00000713;
    mem['h000D] <= 32'h00000793;
    mem['h000E] <= 32'h00000813;
    mem['h000F] <= 32'h00000893;
    mem['h0010] <= 32'h00000913;
    mem['h0011] <= 32'h00000993;
    mem['h0012] <= 32'h00000A13;
    mem['h0013] <= 32'h00000A93;
    mem['h0014] <= 32'h00000B13;
    mem['h0015] <= 32'h00000B93;
    mem['h0016] <= 32'h00000C13;
    mem['h0017] <= 32'h00000C93;
    mem['h0018] <= 32'h00000D13;
    mem['h0019] <= 32'h00000D93;
    mem['h001A] <= 32'h00000E13;
    mem['h001B] <= 32'h00000E93;
    mem['h001C] <= 32'h00000F13;
    mem['h001D] <= 32'h00000F93;
    mem['h001E] <= 32'h00000513;
    mem['h001F] <= 32'h00000593;
    mem['h0020] <= 32'h00B52023;
    mem['h0021] <= 32'h00450513;
    mem['h0022] <= 32'hFE254CE3;
    mem['h0023] <= 32'h00000517;
    mem['h0024] <= 32'h52050513;
    mem['h0025] <= 32'h00000593;
    mem['h0026] <= 32'h01000613;
    mem['h0027] <= 32'h00C5DC63;
    mem['h0028] <= 32'h00052683;
    mem['h0029] <= 32'h00D5A023;
    mem['h002A] <= 32'h00450513;
    mem['h002B] <= 32'h00458593;
    mem['h002C] <= 32'hFEC5C8E3;
    mem['h002D] <= 32'h01000513;
    mem['h002E] <= 32'h01000593;
    mem['h002F] <= 32'h00B55863;
    mem['h0030] <= 32'h00052023;
    mem['h0031] <= 32'h00450513;
    mem['h0032] <= 32'hFEB54CE3;
    mem['h0033] <= 32'h008000EF;
    mem['h0034] <= 32'h0000006F;
    mem['h0035] <= 32'hFF010113;
    mem['h0036] <= 32'h00112623;
    mem['h0037] <= 32'h00812423;
    mem['h0038] <= 32'h01010413;
    mem['h0039] <= 32'h040007B7;
    mem['h003A] <= 32'h01900713;
    mem['h003B] <= 32'h00E7A023;
    mem['h003C] <= 32'h050007B7;
    mem['h003D] <= 32'h01900713;
    mem['h003E] <= 32'h00E7A023;
    mem['h003F] <= 32'h060007B7;
    mem['h0040] <= 32'h06400713;
    mem['h0041] <= 32'h00E7A023;
    mem['h0042] <= 32'h070007B7;
    mem['h0043] <= 32'h06400713;
    mem['h0044] <= 32'h00E7A023;
    mem['h0045] <= 32'h0C0007B7;
    mem['h0046] <= 32'h0007A023;
    mem['h0047] <= 32'h0D0007B7;
    mem['h0048] <= 32'h0007A023;
    mem['h0049] <= 32'h0E0007B7;
    mem['h004A] <= 32'h0007A023;
    mem['h004B] <= 32'h0F0007B7;
    mem['h004C] <= 32'h0007A023;
    mem['h004D] <= 32'h1D8000EF;
    mem['h004E] <= 32'hFFDFF06F;
    mem['h004F] <= 32'hFF010113;
    mem['h0050] <= 32'h00812623;
    mem['h0051] <= 32'h01010413;
    mem['h0052] <= 32'h00802783;
    mem['h0053] <= 32'h01F7D793;
    mem['h0054] <= 32'h0FF7F793;
    mem['h0055] <= 32'h00078513;
    mem['h0056] <= 32'h00C12403;
    mem['h0057] <= 32'h01010113;
    mem['h0058] <= 32'h00008067;
    mem['h0059] <= 32'hFF010113;
    mem['h005A] <= 32'h00812623;
    mem['h005B] <= 32'h01010413;
    mem['h005C] <= 32'h00802783;
    mem['h005D] <= 32'h00F027B3;
    mem['h005E] <= 32'h0FF7F793;
    mem['h005F] <= 32'h00078513;
    mem['h0060] <= 32'h00C12403;
    mem['h0061] <= 32'h01010113;
    mem['h0062] <= 32'h00008067;
    mem['h0063] <= 32'hFF010113;
    mem['h0064] <= 32'h00812623;
    mem['h0065] <= 32'h01010413;
    mem['h0066] <= 32'h060007B7;
    mem['h0067] <= 32'h0007A703;
    mem['h0068] <= 32'h00F00793;
    mem['h0069] <= 32'h02E7EC63;
    mem['h006A] <= 32'h070007B7;
    mem['h006B] <= 32'h0007A703;
    mem['h006C] <= 32'h040007B7;
    mem['h006D] <= 32'h0007A783;
    mem['h006E] <= 32'h02F76263;
    mem['h006F] <= 32'h070007B7;
    mem['h0070] <= 32'h0007A703;
    mem['h0071] <= 32'h040007B7;
    mem['h0072] <= 32'h0007A783;
    mem['h0073] <= 32'h03278793;
    mem['h0074] <= 32'h00E7E663;
    mem['h0075] <= 32'h00100793;
    mem['h0076] <= 32'h0080006F;
    mem['h0077] <= 32'h00000793;
    mem['h0078] <= 32'h0017F793;
    mem['h0079] <= 32'h0FF7F793;
    mem['h007A] <= 32'h00078513;
    mem['h007B] <= 32'h00C12403;
    mem['h007C] <= 32'h01010113;
    mem['h007D] <= 32'h00008067;
    mem['h007E] <= 32'hFF010113;
    mem['h007F] <= 32'h00812623;
    mem['h0080] <= 32'h01010413;
    mem['h0081] <= 32'h060007B7;
    mem['h0082] <= 32'h0007A703;
    mem['h0083] <= 32'h26600793;
    mem['h0084] <= 32'h02E7FC63;
    mem['h0085] <= 32'h070007B7;
    mem['h0086] <= 32'h0007A703;
    mem['h0087] <= 32'h050007B7;
    mem['h0088] <= 32'h0007A783;
    mem['h0089] <= 32'h02F76263;
    mem['h008A] <= 32'h070007B7;
    mem['h008B] <= 32'h0007A703;
    mem['h008C] <= 32'h050007B7;
    mem['h008D] <= 32'h0007A783;
    mem['h008E] <= 32'h03278793;
    mem['h008F] <= 32'h00E7E663;
    mem['h0090] <= 32'h00100793;
    mem['h0091] <= 32'h0080006F;
    mem['h0092] <= 32'h00000793;
    mem['h0093] <= 32'h0017F793;
    mem['h0094] <= 32'h0FF7F793;
    mem['h0095] <= 32'h00078513;
    mem['h0096] <= 32'h00C12403;
    mem['h0097] <= 32'h01010113;
    mem['h0098] <= 32'h00008067;
    mem['h0099] <= 32'hFF010113;
    mem['h009A] <= 32'h00812623;
    mem['h009B] <= 32'h01010413;
    mem['h009C] <= 32'h0D0007B7;
    mem['h009D] <= 32'h0007A703;
    mem['h009E] <= 32'h00170713;
    mem['h009F] <= 32'h00E7A023;
    mem['h00A0] <= 32'h0D0007B7;
    mem['h00A1] <= 32'h0007A703;
    mem['h00A2] <= 32'h00900793;
    mem['h00A3] <= 32'h00E7FE63;
    mem['h00A4] <= 32'h0D0007B7;
    mem['h00A5] <= 32'h0007A023;
    mem['h00A6] <= 32'h0C0007B7;
    mem['h00A7] <= 32'h0007A703;
    mem['h00A8] <= 32'h00170713;
    mem['h00A9] <= 32'h00E7A023;
    mem['h00AA] <= 32'h00000013;
    mem['h00AB] <= 32'h00C12403;
    mem['h00AC] <= 32'h01010113;
    mem['h00AD] <= 32'h00008067;
    mem['h00AE] <= 32'hFF010113;
    mem['h00AF] <= 32'h00812623;
    mem['h00B0] <= 32'h01010413;
    mem['h00B1] <= 32'h0F0007B7;
    mem['h00B2] <= 32'h0007A703;
    mem['h00B3] <= 32'h00170713;
    mem['h00B4] <= 32'h00E7A023;
    mem['h00B5] <= 32'h0F0007B7;
    mem['h00B6] <= 32'h0007A703;
    mem['h00B7] <= 32'h00900793;
    mem['h00B8] <= 32'h00E7FE63;
    mem['h00B9] <= 32'h0F0007B7;
    mem['h00BA] <= 32'h0007A023;
    mem['h00BB] <= 32'h0E0007B7;
    mem['h00BC] <= 32'h0007A703;
    mem['h00BD] <= 32'h00170713;
    mem['h00BE] <= 32'h00E7A023;
    mem['h00BF] <= 32'h00000013;
    mem['h00C0] <= 32'h00C12403;
    mem['h00C1] <= 32'h01010113;
    mem['h00C2] <= 32'h00008067;
    mem['h00C3] <= 32'hFF010113;
    mem['h00C4] <= 32'h00112623;
    mem['h00C5] <= 32'h00812423;
    mem['h00C6] <= 32'h01010413;
    mem['h00C7] <= 32'h00002783;
    mem['h00C8] <= 32'hFFF78713;
    mem['h00C9] <= 32'h00E02023;
    mem['h00CA] <= 32'h00402783;
    mem['h00CB] <= 32'hFFF78713;
    mem['h00CC] <= 32'h00E02223;
    mem['h00CD] <= 32'h00402783;
    mem['h00CE] <= 32'h04079463;
    mem['h00CF] <= 32'h00001737;
    mem['h00D0] <= 32'h77070713;
    mem['h00D1] <= 32'h00E02223;
    mem['h00D2] <= 32'h060007B7;
    mem['h00D3] <= 32'h0007A703;
    mem['h00D4] <= 32'h00802783;
    mem['h00D5] <= 32'h00078693;
    mem['h00D6] <= 32'h060007B7;
    mem['h00D7] <= 32'h00D70733;
    mem['h00D8] <= 32'h00E7A023;
    mem['h00D9] <= 32'h070007B7;
    mem['h00DA] <= 32'h0007A703;
    mem['h00DB] <= 32'h00C02783;
    mem['h00DC] <= 32'h00078693;
    mem['h00DD] <= 32'h070007B7;
    mem['h00DE] <= 32'h00D70733;
    mem['h00DF] <= 32'h00E7A023;
    mem['h00E0] <= 32'h00002783;
    mem['h00E1] <= 32'h20079A63;
    mem['h00E2] <= 32'h00001737;
    mem['h00E3] <= 32'hFA070713;
    mem['h00E4] <= 32'h00E02023;
    mem['h00E5] <= 32'h0C0007B7;
    mem['h00E6] <= 32'h0007A703;
    mem['h00E7] <= 32'h00900793;
    mem['h00E8] <= 32'h02F71A63;
    mem['h00E9] <= 32'h0D0007B7;
    mem['h00EA] <= 32'h0007A703;
    mem['h00EB] <= 32'h00900793;
    mem['h00EC] <= 32'h02F71263;
    mem['h00ED] <= 32'h0C0007B7;
    mem['h00EE] <= 32'h0007A023;
    mem['h00EF] <= 32'h0D0007B7;
    mem['h00F0] <= 32'h0007A023;
    mem['h00F1] <= 32'h0E0007B7;
    mem['h00F2] <= 32'h0007A023;
    mem['h00F3] <= 32'h0F0007B7;
    mem['h00F4] <= 32'h0007A023;
    mem['h00F5] <= 32'h0E0007B7;
    mem['h00F6] <= 32'h0007A703;
    mem['h00F7] <= 32'h00900793;
    mem['h00F8] <= 32'h02F71A63;
    mem['h00F9] <= 32'h0F0007B7;
    mem['h00FA] <= 32'h0007A703;
    mem['h00FB] <= 32'h00900793;
    mem['h00FC] <= 32'h02F71263;
    mem['h00FD] <= 32'h0C0007B7;
    mem['h00FE] <= 32'h0007A023;
    mem['h00FF] <= 32'h0D0007B7;
    mem['h0100] <= 32'h0007A023;
    mem['h0101] <= 32'h0E0007B7;
    mem['h0102] <= 32'h0007A023;
    mem['h0103] <= 32'h0F0007B7;
    mem['h0104] <= 32'h0007A023;
    mem['h0105] <= 32'h080007B7;
    mem['h0106] <= 32'h0007A703;
    mem['h0107] <= 32'h00100793;
    mem['h0108] <= 32'h02F71063;
    mem['h0109] <= 32'h040007B7;
    mem['h010A] <= 32'h0007A783;
    mem['h010B] <= 32'h00078A63;
    mem['h010C] <= 32'h040007B7;
    mem['h010D] <= 32'h0007A703;
    mem['h010E] <= 32'hFFF70713;
    mem['h010F] <= 32'h00E7A023;
    mem['h0110] <= 32'h090007B7;
    mem['h0111] <= 32'h0007A703;
    mem['h0112] <= 32'h00100793;
    mem['h0113] <= 32'h02F71263;
    mem['h0114] <= 32'h040007B7;
    mem['h0115] <= 32'h0007A703;
    mem['h0116] <= 32'h1AD00793;
    mem['h0117] <= 32'h00E7EA63;
    mem['h0118] <= 32'h040007B7;
    mem['h0119] <= 32'h0007A703;
    mem['h011A] <= 32'h00170713;
    mem['h011B] <= 32'h00E7A023;
    mem['h011C] <= 32'h0A0007B7;
    mem['h011D] <= 32'h0007A703;
    mem['h011E] <= 32'h00100793;
    mem['h011F] <= 32'h02F71063;
    mem['h0120] <= 32'h050007B7;
    mem['h0121] <= 32'h0007A783;
    mem['h0122] <= 32'h00078A63;
    mem['h0123] <= 32'h050007B7;
    mem['h0124] <= 32'h0007A703;
    mem['h0125] <= 32'hFFF70713;
    mem['h0126] <= 32'h00E7A023;
    mem['h0127] <= 32'h0B0007B7;
    mem['h0128] <= 32'h0007A703;
    mem['h0129] <= 32'h00100793;
    mem['h012A] <= 32'h02F71263;
    mem['h012B] <= 32'h050007B7;
    mem['h012C] <= 32'h0007A703;
    mem['h012D] <= 32'h1AD00793;
    mem['h012E] <= 32'h00E7EA63;
    mem['h012F] <= 32'h050007B7;
    mem['h0130] <= 32'h0007A703;
    mem['h0131] <= 32'h00170713;
    mem['h0132] <= 32'h00E7A023;
    mem['h0133] <= 32'h070007B7;
    mem['h0134] <= 32'h0007A703;
    mem['h0135] <= 32'h01900793;
    mem['h0136] <= 32'h00E7FA63;
    mem['h0137] <= 32'h070007B7;
    mem['h0138] <= 32'h0007A703;
    mem['h0139] <= 32'h1DF00793;
    mem['h013A] <= 32'h00E7F863;
    mem['h013B] <= 32'h00C02783;
    mem['h013C] <= 32'h40F00733;
    mem['h013D] <= 32'h00E02623;
    mem['h013E] <= 32'hC45FF0EF;
    mem['h013F] <= 32'h00050793;
    mem['h0140] <= 32'h00078E63;
    mem['h0141] <= 32'hC89FF0EF;
    mem['h0142] <= 32'h00050793;
    mem['h0143] <= 32'h00078863;
    mem['h0144] <= 32'h00802783;
    mem['h0145] <= 32'h40F00733;
    mem['h0146] <= 32'h00E02423;
    mem['h0147] <= 32'hC49FF0EF;
    mem['h0148] <= 32'h00050793;
    mem['h0149] <= 32'h00078E63;
    mem['h014A] <= 32'hCD1FF0EF;
    mem['h014B] <= 32'h00050793;
    mem['h014C] <= 32'h00078863;
    mem['h014D] <= 32'h00802783;
    mem['h014E] <= 32'h40F00733;
    mem['h014F] <= 32'h00E02423;
    mem['h0150] <= 32'h060007B7;
    mem['h0151] <= 32'h0007A783;
    mem['h0152] <= 32'h00078A63;
    mem['h0153] <= 32'h060007B7;
    mem['h0154] <= 32'h0007A703;
    mem['h0155] <= 32'h27F00793;
    mem['h0156] <= 32'h04E7F063;
    mem['h0157] <= 32'hBE1FF0EF;
    mem['h0158] <= 32'h00050793;
    mem['h0159] <= 32'h00078663;
    mem['h015A] <= 32'hD51FF0EF;
    mem['h015B] <= 32'h0080006F;
    mem['h015C] <= 32'hCF5FF0EF;
    mem['h015D] <= 32'h00802783;
    mem['h015E] <= 32'h40F00733;
    mem['h015F] <= 32'h00E02423;
    mem['h0160] <= 32'h060007B7;
    mem['h0161] <= 32'h14000713;
    mem['h0162] <= 32'h00E7A023;
    mem['h0163] <= 32'h070007B7;
    mem['h0164] <= 32'h0F000713;
    mem['h0165] <= 32'h00E7A023;
    mem['h0166] <= 32'h00000013;
    mem['h0167] <= 32'h00C12083;
    mem['h0168] <= 32'h00812403;
    mem['h0169] <= 32'h01010113;
    mem['h016A] <= 32'h00008067;
    mem['h016B] <= 32'h00000FA0;
    mem['h016C] <= 32'h00001770;
    mem['h016D] <= 32'h00000001;
    mem['h016E] <= 32'h00000001;

  end

  always @(posedge clk) mem_data <= mem[mem_addr];

  // ============================================================================

  reg o_ready;

  always @(posedge clk or negedge rstn)
    if (!rstn) o_ready <= 1'd0;
    else o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

  // Output connectins
  assign ready    = o_ready;
  assign rdata    = mem_data;
  assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule
